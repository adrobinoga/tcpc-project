module tcpc();

//------------------------------------------------------------
// Registros

wire [15:0] RD_DATA;
wire [15:0] WR_DATA;
wire [7:0] ADDR;
wire [15:0] DEVICE_ID;
wire [15:0] USBTYPEC_REV;
wire [15:0] USBPD_REV_VER;
wire [15:0] PD_INTERFACE_REV;
wire [15:0] ALERT;
wire [15:0] ALERT_MASK;
wire [7:0] POWER_STATUS_MASK;
wire [7:0] FAULT_STATUS_MASK;
output [7:0] TCPC_CONTROL;
wire [7:0] ROLE_CONTROL;
wire [7:0] FAULT_CONTROL;
wire [7:0] POWER_CONTROL;
wire [7:0] CC_STATUS;
wire [7:0] POWER_STATUS;
wire [7:0] FAULT_STATUS;
wire [15:0] Reserved;
wire [7:0] COMMAND;
wire [15:0] DEVICE_CAPABILITIES_1;
wire [15:0] DEVICE_CAPABILITIES_2;
wire [7:0] STANDARD_INPUT_CAPABILITIES;
wire [15:0] STANDARD_OUTPUT_CAPABILITIES;
wire [7:0] MESSAGE_HEADER_INFO;
wire [7:0] RECEIVE_DETECT;
wire [7:0] RECEIVE_BYTE_COUNT;
wire [7:0] RX_BUF_FRAME_TYPE;
wire [7:0] RX_BUF_HEADER_BYTE_0;
wire [7:0] RX_BUF_HEADER_BYTE_1;
wire [7:0] RX_BUF_OBJ1_BYTE_0;
wire [7:0] RX_BUF_OBJ1_BYTE_1;
wire [7:0] RX_BUF_OBJ1_BYTE_2;
wire [7:0] RX_BUF_OBJ1_BYTE_3;
wire [7:0] RX_BUF_OBJ2_BYTE_0;
wire [15:0] RX_BUF_OBJn_BYTE_m;
wire [7:0] RX_BUF_OBJ7_BYTE_3;
wire [7:0] TRANSMIT;
wire [7:0] TRANSMIT_BYTE_COUNT;
wire [7:0] TX_BUF_HEADER_BYTE_0;	
wire [7:0] TX_BUF_HEADER_BYTE_1;
wire [7:0] TX_BUF_OBJ1_BYTE_0;
wire [15:0] TX_BUF_OBJn_BYTE_m;
wire [7:0] TX_BUF_OBJ7_BYTE_3;
wire [15:0] VBUS_VOLTAGE;
wire [15:0] VBUS_SINK_DISCONNECT_THRESHOLD;
wire [15:0] VBUS_STOP_DISCHARGE_THRESHOLD;
wire [15:0] VBUS_SINK_DISCHARGE_THRESHOLD;
wire [15:0] VBUS_VOLTAGE_ALARM_HI_CFG;
wire [15:0] VBUS_VOLTAGE_ALARM_LO_CFG;
//------------------------------------------------------------

rx rxu();

tx txu();

i2c_slave i2c_slave_u();

registers registers_u(
	.CLK(CLK),
	.RNW(RNW), 
	.WR_DATA(WR_DATA),
	.RD_DATA(RD_DATA), 
	.REQUEST(REQUEST), 
	.ADDR(ADDR),
	.ACK(ACK),
	
	// registros de uso inmediato
	.DEVICE_ID(DEVICE_ID),      				              		
	.USBTYPEC_REV(USBTYPEC_REV),					    	
	.USBPD_REV_VER(USBPD_REV_VER),				    		
	.PD_INTERFACE_REV(PD_INTERFACE_REV),			   		
	.ALERT(ALERT),						    		
	.ALERT_MASK(ALERT_MASK),				    		
	.POWER_STATUS_MASK(POWER_STATUS_MASK),			    	
	.FAULT_STATUS_MASK(FAULT_STATUS_MASK),			    	  		
	.TCPC_CONTROL(TCPC_CONTROL),				    		
	.ROLE_CONTROL(ROLE_CONTROL),				    		
	.FAULT_CONTROL(FAULT_CONTROL),				    		
	.POWER_CONTROL(POWER_CONTROL),				    		
	.CC_STATUS(CC_STATUS),					    		
	.POWER_STATUS(POWER_STATUS),				    		
	.FAULT_STATUS(FAULT_STATUS),					 		    
	.COMMAND(COMMAND),							    	
	.DEVICE_CAPABILITIES_1(DEVICE_CAPABILITIES_1), 		 	  		
	.DEVICE_CAPABILITIES_2(DEVICE_CAPABILITIES_2), 		   		
	.STANDARD_INPUT_CAPABILITIES(STANDARD_INPUT_CAPABILITIES), 	  	
	.STANDARD_OUTPUT_CAPABILITIES(STANDARD_OUTPUT_CAPABILITIES), 	  		
	.MESSAGE_HEADER_INFO(MESSAGE_HEADER_INFO), 					
	.RECEIVE_DETECT(RECEIVE_DETECT), 						
	.RECEIVE_BYTE_COUNT(RECEIVE_BYTE_COUNT), 			 		

	.RX_BUF_FRAME_TYPE(RX_BUF_FRAME_TYPE), 					
	.RX_BUF_HEADER_BYTE_0(RX_BUF_HEADER_BYTE_0), 			 		
	.RX_BUF_HEADER_BYTE_1(RX_BUF_HEADER_BYTE_1),			  	
	.RX_BUF_OBJ1_BYTE_0(RX_BUF_OBJ1_BYTE_0), 			 		
	.RX_BUF_OBJ1_BYTE_1(RX_BUF_OBJ1_BYTE_1),			  		
	.RX_BUF_OBJ1_BYTE_2(RX_BUF_OBJ1_BYTE_2), 			 		
	.RX_BUF_OBJ1_BYTE_3(RX_BUF_OBJ1_BYTE_3),			 	
	.RX_BUF_OBJ2_BYTE_0(RX_BUF_OBJ2_BYTE_0),			 	
	.RX_BUF_OBJ2_BYTE_1(RX_BUF_OBJ2_BYTE_1),			 	
	.RX_BUF_OBJ2_BYTE_2(RX_BUF_OBJ2_BYTE_2),			 	
	.RX_BUF_OBJ2_BYTE_3(RX_BUF_OBJ2_BYTE_3), 			 		

	.TRANSMIT(TRANSMIT),							
	.TRANSMIT_BYTE_COUNT(TRANSMIT_BYTE_COUNT), 	
				
	.TX_BUF_HEADER_BYTE_0(TX_BUF_HEADER_BYTE_0), 			
	.TX_BUF_HEADER_BYTE_1(TX_BUF_HEADER_BYTE_1), 	
	.TX_BUF_OBJ1_BYTE_0(TX_BUF_OBJ1_BYTE_0), 			 		
	.TX_BUF_OBJ1_BYTE_1(TX_BUF_OBJ1_BYTE_1),			  		
	.TX_BUF_OBJ1_BYTE_2(TX_BUF_OBJ1_BYTE_2), 			 		
	.TX_BUF_OBJ1_BYTE_3(TX_BUF_OBJ1_BYTE_3),			 	
	.TX_BUF_OBJ2_BYTE_0(TX_BUF_OBJ2_BYTE_0),			 	
	.TX_BUF_OBJ2_BYTE_1(TX_BUF_OBJ2_BYTE_1),			 	
	.TX_BUF_OBJ2_BYTE_2(TX_BUF_OBJ2_BYTE_2),			 	
	.TX_BUF_OBJ2_BYTE_3(TX_BUF_OBJ2_BYTE_3),					
	
	.VBUS_VOLTAGE(VBUS_VOLTAGE)
	); 	

endmodule
