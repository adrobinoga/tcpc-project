
module tester(
	
);

initial
	begin
	
	
	end
endmodule
