module tcpc();

rx rxu();

tx txu();

i2c_slave i2c_slave_u();

registers registers_u();

endmodule
